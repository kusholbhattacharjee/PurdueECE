// $Id: $
// File name:   tb_usb_receiver.sv
// Created:     2/28/2018
// Author:      Kushol Bhattacharjee
// Lab Section: 337-07
// Version:     1.0  Initial Design Entry
// Description: test bench for usb_receiver.sv

`timescale 1ns/ 100 ps 

module tb_usb_receiver(); 

endmodule 
