// $Id: $
// File name:   tb_rx_fifo.sv
// Created:     2/21/2018
// Author:      Kushol Bhattacharjee
// Lab Section: 337-07
// Version:     1.0  Initial Design Entry
// Description: top level test bench for rx_fifo

`timescale 1ns/ 100 ps

module tb_rx_fifo(); 

endmodule
